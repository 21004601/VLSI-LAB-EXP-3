module multiplier_4bit(
input [3:0] a, b,
output [7:0] result
);
assign result = a * b;
endmodule





